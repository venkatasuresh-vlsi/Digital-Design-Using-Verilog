module comp (
     input a, b,
	 output eq
	 );
	 xnor G4 (eq, a, b);
	 
	endmodule