module tb;
     reg clk, rst, inc;
	 reg [2:0] val;
	 wire [7:0] cnt;
	 reg incNBA;
	 
	 always @* incNBA <=inc;
	 
	 inc_by_value Suresh (clk, rst, incNBA, val, cnt);
	 
	 always #5 clk = !clk;
	 initial clk = 0;
	 
	 initial begin
	     rst = 1; inc = 0; val = 2'b00; #10;
		 rst = 0;
		 @(posedge clk);
		 @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd3; @(negedge clk); inc = 0; val = 3'd3; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd4; @(negedge clk); inc = 0; val = 3'd4; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd5; @(negedge clk); inc = 0; val = 3'd5; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd6; @(negedge clk); inc = 0; val = 3'd6; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd7; @(negedge clk); inc = 0; val = 3'd7; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd1; @(negedge clk); inc = 0; val = 3'd1; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd2; @(negedge clk); inc = 0; val = 3'd3; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd4; @(negedge clk); inc = 0; val = 3'd3; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd5; @(negedge clk); inc = 0; val = 3'd3; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd6; @(negedge clk); inc = 0; val = 3'd3; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd5; @(negedge clk); inc = 0; val = 3'd3; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd4; @(negedge clk); inc = 0; val = 3'd3; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd3; @(negedge clk); inc = 0; val = 3'd3; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd2; @(negedge clk); inc = 0; val = 3'd3; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd1; @(negedge clk); inc = 0; val = 3'd3; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd0; @(negedge clk); inc = 0; val = 3'd3; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd2; @(negedge clk); inc = 0; val = 3'd3; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd7; @(negedge clk); inc = 0; val = 3'd3; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd6; @(negedge clk); inc = 0; val = 3'd3; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd4; @(negedge clk); inc = 0; val = 3'd5; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd5; @(negedge clk); inc = 0; val = 3'd5; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd6; @(negedge clk); inc = 0; val = 3'd4; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd2; @(negedge clk); inc = 0; val = 3'd3; 
         @(posedge clk);
		 @(posedge clk);
		 @(negedge clk); inc = 1; val = 3'd0; @(negedge clk); inc = 0; val = 3'd0; 
         @(posedge clk);
		 @(posedge clk);
		 $finish;
		end
	endmodule